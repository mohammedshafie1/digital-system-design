LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_arith.all;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY ASSIGNMENT IS
PORT(
		X,Y      :IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		SEG1,SEG2:BUFFER STD_LOGIC_VECTOR(0 TO 6);
		F : BUFFER STD_LOGIC_VECTOR(4 DOWNTO 0)
    );
END ASSIGNMENT;



ARCHITECTURE ASSIGNMENT_ARCH OF ASSIGNMENT IS
SIGNAL Z: STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL S:STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL S1:STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL S2:STD_LOGIC_VECTOR(3 DOWNTO 0);

BEGIN

 PROCESS(X,Y)
 BEGIN
   
	Z<=('0' & X) + Y;
	F<=Z;
	
	

	CASE F IS
	 WHEN "00000" => SEG1 <="0000001";SEG2<="0000001";
	 WHEN "00001" => SEG1 <="1001111";SEG2<="0000001";
	 WHEN "00010" => SEG1 <="0010010";SEG2<="0000001";
	 WHEN "00011" => SEG1 <="0000110";SEG2<="0000001";
	 WHEN "00100" => SEG1 <="1001100";SEG2<="0000001";
	 WHEN "00101" => SEG1 <="0100100";SEG2<="0000001";
	 WHEN "00110" => SEG1 <="0100000";SEG2<="0000001";
	 WHEN "00111" => SEG1 <="0001111";SEG2<="0000001";
	 WHEN "01000" => SEG1 <="0000000";SEG2<="0000001";
	 WHEN "01001" => SEG1 <="0000100";SEG2<="0000001";
	 
	 
	 
	 WHEN "01010" => SEG1 <="0000001";SEG2<="1001111";
	 WHEN "01011" => SEG1 <="1001111";SEG2<="1001111";
	 WHEN "01100" => SEG1 <="0010010";SEG2<="1001111";
	 WHEN "01101" => SEG1 <="0000110";SEG2<="1001111";
	 WHEN "01110" => SEG1 <="1001100";SEG2<="1001111";
	 WHEN "01111" => SEG1 <="0100100";SEG2<="1001111";
	 WHEN "10000" => SEG1 <="0100000";SEG2<="1001111";
	 WHEN "10001" => SEG1 <="0001111";SEG2<="1001111";
	 WHEN "10010" => SEG1 <="0000000";SEG2<="1001111";
	 WHEN "10011" => SEG1 <="0000100";SEG2<="1001111";
	 
	 
	 WHEN "10100" => SEG1 <="0000001";SEG2<="0010010";
	 WHEN "10101" => SEG1 <="1001111";SEG2<="0010010";
	 WHEN "10110" => SEG1 <="0010010";SEG2<="0010010";
	 WHEN "10111" => SEG1 <="0000110";SEG2<="0010010";
	 WHEN "11000" => SEG1 <="1001100";SEG2<="0010010";
	 WHEN "11001" => SEG1 <="0100100";SEG2<="0010010";
	 WHEN "11010" => SEG1 <="0100000";SEG2<="0010010";
	 WHEN "11011" => SEG1 <="0001111";SEG2<="0010010";
	 WHEN "11100" => SEG1 <="0000000";SEG2<="0010010";
	 WHEN "11101" => SEG1 <="0000100";SEG2<="0010010";
	 
	 WHEN "11110" => SEG1 <="0000001";SEG2<="0000110";
	 WHEN OTHERS => SEG1 <= "-------";SEG2<="-------";
	
	 
 END CASE;	
 END PROCESS;

END ASSIGNMENT_ARCH;